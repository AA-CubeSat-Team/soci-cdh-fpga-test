
module NIOS_2 (
	clk_clk);	

	input		clk_clk;
endmodule
