module NIOS_2_Top (
	input  		MAX10_CLK1_50
);
	NIOS_2 nios (.clk_clk(MAX10_CLK1_50));
endmodule 